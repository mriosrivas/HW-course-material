//HDL Example 4.26 PRIORITY CIRCUIT

module priorityckt(input logic [3:0] a,
    output logic [3:0] y);

    always_comb
        if      (a[3]) y <= 4'b1000;
        else if (a[2]) y <= 4'b0100;
        else if (a[1]) y <= 4'b0010;
        else if (a[0]) y <= 4'b0001;
        else y <= 4'b0000;
        
endmodule